magic
tech scmos
timestamp 1619554542
<< nwell >>
rect -341 292 -243 324
rect -205 297 -107 329
rect -341 184 -287 216
rect -223 177 -169 209
rect -96 199 2 231
rect -341 114 -243 146
rect -160 106 -106 138
rect -92 42 -38 74
rect -341 6 -287 38
rect 35 27 133 59
rect -29 -17 25 15
rect -341 -64 -243 -32
rect 40 -81 94 -49
rect 109 -138 163 -106
rect -341 -172 -287 -140
rect -341 -242 -243 -210
rect -341 -350 -287 -318
<< ntransistor >>
rect -329 275 -327 285
rect -257 275 -255 285
rect -193 280 -191 290
rect -121 280 -119 290
rect -305 240 -303 250
rect -295 240 -293 250
rect -285 240 -283 250
rect -275 240 -273 250
rect -169 245 -167 255
rect -159 245 -157 255
rect -149 245 -147 255
rect -139 245 -137 255
rect -329 160 -327 170
rect -319 160 -317 170
rect -301 160 -299 170
rect -84 182 -82 192
rect -211 153 -209 163
rect -201 153 -199 163
rect -183 153 -181 163
rect -12 182 -10 192
rect -60 147 -58 157
rect -50 147 -48 157
rect -40 147 -38 157
rect -30 147 -28 157
rect -329 97 -327 107
rect -257 97 -255 107
rect -148 82 -146 92
rect -138 82 -136 92
rect -120 82 -118 92
rect -305 62 -303 72
rect -295 62 -293 72
rect -285 62 -283 72
rect -275 62 -273 72
rect -80 18 -78 28
rect -70 18 -68 28
rect -52 18 -50 28
rect 47 10 49 20
rect -329 -18 -327 -8
rect -319 -18 -317 -8
rect -301 -18 -299 -8
rect 119 10 121 20
rect 71 -25 73 -15
rect 81 -25 83 -15
rect 91 -25 93 -15
rect 101 -25 103 -15
rect -17 -41 -15 -31
rect -7 -41 -5 -31
rect 11 -41 13 -31
rect -329 -81 -327 -71
rect -257 -81 -255 -71
rect 52 -105 54 -95
rect 62 -105 64 -95
rect 80 -105 82 -95
rect -305 -116 -303 -106
rect -295 -116 -293 -106
rect -285 -116 -283 -106
rect -275 -116 -273 -106
rect 121 -162 123 -152
rect 131 -162 133 -152
rect 149 -162 151 -152
rect -329 -196 -327 -186
rect -319 -196 -317 -186
rect -301 -196 -299 -186
rect -329 -259 -327 -249
rect -257 -259 -255 -249
rect -305 -294 -303 -284
rect -295 -294 -293 -284
rect -285 -294 -283 -284
rect -275 -294 -273 -284
rect -329 -374 -327 -364
rect -319 -374 -317 -364
rect -301 -374 -299 -364
<< ptransistor >>
rect -329 298 -327 318
rect -305 298 -303 318
rect -295 298 -293 318
rect -285 298 -283 318
rect -275 298 -273 318
rect -257 298 -255 318
rect -193 303 -191 323
rect -169 303 -167 323
rect -159 303 -157 323
rect -149 303 -147 323
rect -139 303 -137 323
rect -121 303 -119 323
rect -329 190 -327 210
rect -319 190 -317 210
rect -301 190 -299 210
rect -84 205 -82 225
rect -60 205 -58 225
rect -50 205 -48 225
rect -40 205 -38 225
rect -30 205 -28 225
rect -12 205 -10 225
rect -211 183 -209 203
rect -201 183 -199 203
rect -183 183 -181 203
rect -329 120 -327 140
rect -305 120 -303 140
rect -295 120 -293 140
rect -285 120 -283 140
rect -275 120 -273 140
rect -257 120 -255 140
rect -148 112 -146 132
rect -138 112 -136 132
rect -120 112 -118 132
rect -80 48 -78 68
rect -70 48 -68 68
rect -52 48 -50 68
rect -329 12 -327 32
rect -319 12 -317 32
rect -301 12 -299 32
rect 47 33 49 53
rect 71 33 73 53
rect 81 33 83 53
rect 91 33 93 53
rect 101 33 103 53
rect 119 33 121 53
rect -17 -11 -15 9
rect -7 -11 -5 9
rect 11 -11 13 9
rect -329 -58 -327 -38
rect -305 -58 -303 -38
rect -295 -58 -293 -38
rect -285 -58 -283 -38
rect -275 -58 -273 -38
rect -257 -58 -255 -38
rect 52 -75 54 -55
rect 62 -75 64 -55
rect 80 -75 82 -55
rect 121 -132 123 -112
rect 131 -132 133 -112
rect 149 -132 151 -112
rect -329 -166 -327 -146
rect -319 -166 -317 -146
rect -301 -166 -299 -146
rect -329 -236 -327 -216
rect -305 -236 -303 -216
rect -295 -236 -293 -216
rect -285 -236 -283 -216
rect -275 -236 -273 -216
rect -257 -236 -255 -216
rect -329 -344 -327 -324
rect -319 -344 -317 -324
rect -301 -344 -299 -324
<< ndiffusion >>
rect -331 275 -329 285
rect -327 275 -325 285
rect -259 275 -257 285
rect -255 275 -253 285
rect -195 280 -193 290
rect -191 280 -189 290
rect -123 280 -121 290
rect -119 280 -117 290
rect -307 240 -305 250
rect -303 240 -301 250
rect -297 240 -295 250
rect -293 240 -291 250
rect -287 240 -285 250
rect -283 240 -281 250
rect -277 240 -275 250
rect -273 240 -271 250
rect -171 245 -169 255
rect -167 245 -165 255
rect -161 245 -159 255
rect -157 245 -155 255
rect -151 245 -149 255
rect -147 245 -145 255
rect -141 245 -139 255
rect -137 245 -135 255
rect -331 160 -329 170
rect -327 160 -319 170
rect -317 160 -315 170
rect -303 160 -301 170
rect -299 160 -297 170
rect -86 182 -84 192
rect -82 182 -80 192
rect -213 153 -211 163
rect -209 153 -201 163
rect -199 153 -197 163
rect -185 153 -183 163
rect -181 153 -179 163
rect -14 182 -12 192
rect -10 182 -8 192
rect -62 147 -60 157
rect -58 147 -56 157
rect -52 147 -50 157
rect -48 147 -46 157
rect -42 147 -40 157
rect -38 147 -36 157
rect -32 147 -30 157
rect -28 147 -26 157
rect -331 97 -329 107
rect -327 97 -325 107
rect -259 97 -257 107
rect -255 97 -253 107
rect -150 82 -148 92
rect -146 82 -144 92
rect -140 82 -138 92
rect -136 82 -134 92
rect -122 82 -120 92
rect -118 82 -116 92
rect -307 62 -305 72
rect -303 62 -301 72
rect -297 62 -295 72
rect -293 62 -291 72
rect -287 62 -285 72
rect -283 62 -281 72
rect -277 62 -275 72
rect -273 62 -271 72
rect -82 18 -80 28
rect -78 18 -70 28
rect -68 18 -66 28
rect -54 18 -52 28
rect -50 18 -48 28
rect 45 10 47 20
rect 49 10 51 20
rect -331 -18 -329 -8
rect -327 -18 -319 -8
rect -317 -18 -315 -8
rect -303 -18 -301 -8
rect -299 -18 -297 -8
rect 117 10 119 20
rect 121 10 123 20
rect 69 -25 71 -15
rect 73 -25 75 -15
rect 79 -25 81 -15
rect 83 -25 85 -15
rect 89 -25 91 -15
rect 93 -25 95 -15
rect 99 -25 101 -15
rect 103 -25 105 -15
rect -19 -41 -17 -31
rect -15 -41 -13 -31
rect -9 -41 -7 -31
rect -5 -41 -3 -31
rect 9 -41 11 -31
rect 13 -41 15 -31
rect -331 -81 -329 -71
rect -327 -81 -325 -71
rect -259 -81 -257 -71
rect -255 -81 -253 -71
rect 50 -105 52 -95
rect 54 -105 62 -95
rect 64 -105 66 -95
rect 78 -105 80 -95
rect 82 -105 84 -95
rect -307 -116 -305 -106
rect -303 -116 -301 -106
rect -297 -116 -295 -106
rect -293 -116 -291 -106
rect -287 -116 -285 -106
rect -283 -116 -281 -106
rect -277 -116 -275 -106
rect -273 -116 -271 -106
rect 119 -162 121 -152
rect 123 -162 125 -152
rect 129 -162 131 -152
rect 133 -162 135 -152
rect 147 -162 149 -152
rect 151 -162 153 -152
rect -331 -196 -329 -186
rect -327 -196 -319 -186
rect -317 -196 -315 -186
rect -303 -196 -301 -186
rect -299 -196 -297 -186
rect -331 -259 -329 -249
rect -327 -259 -325 -249
rect -259 -259 -257 -249
rect -255 -259 -253 -249
rect -307 -294 -305 -284
rect -303 -294 -301 -284
rect -297 -294 -295 -284
rect -293 -294 -291 -284
rect -287 -294 -285 -284
rect -283 -294 -281 -284
rect -277 -294 -275 -284
rect -273 -294 -271 -284
rect -331 -374 -329 -364
rect -327 -374 -319 -364
rect -317 -374 -315 -364
rect -303 -374 -301 -364
rect -299 -374 -297 -364
<< pdiffusion >>
rect -331 298 -329 318
rect -327 298 -325 318
rect -307 298 -305 318
rect -303 298 -295 318
rect -293 298 -291 318
rect -287 298 -285 318
rect -283 298 -275 318
rect -273 298 -271 318
rect -259 298 -257 318
rect -255 298 -253 318
rect -195 303 -193 323
rect -191 303 -189 323
rect -171 303 -169 323
rect -167 303 -159 323
rect -157 303 -155 323
rect -151 303 -149 323
rect -147 303 -139 323
rect -137 303 -135 323
rect -123 303 -121 323
rect -119 303 -117 323
rect -331 190 -329 210
rect -327 190 -325 210
rect -321 190 -319 210
rect -317 190 -315 210
rect -303 190 -301 210
rect -299 190 -297 210
rect -86 205 -84 225
rect -82 205 -80 225
rect -62 205 -60 225
rect -58 205 -50 225
rect -48 205 -46 225
rect -42 205 -40 225
rect -38 205 -30 225
rect -28 205 -26 225
rect -14 205 -12 225
rect -10 205 -8 225
rect -213 183 -211 203
rect -209 183 -207 203
rect -203 183 -201 203
rect -199 183 -197 203
rect -185 183 -183 203
rect -181 183 -179 203
rect -331 120 -329 140
rect -327 120 -325 140
rect -307 120 -305 140
rect -303 120 -295 140
rect -293 120 -291 140
rect -287 120 -285 140
rect -283 120 -275 140
rect -273 120 -271 140
rect -259 120 -257 140
rect -255 120 -253 140
rect -150 112 -148 132
rect -146 112 -138 132
rect -136 112 -134 132
rect -122 112 -120 132
rect -118 112 -116 132
rect -82 48 -80 68
rect -78 48 -76 68
rect -72 48 -70 68
rect -68 48 -66 68
rect -54 48 -52 68
rect -50 48 -48 68
rect -331 12 -329 32
rect -327 12 -325 32
rect -321 12 -319 32
rect -317 12 -315 32
rect -303 12 -301 32
rect -299 12 -297 32
rect 45 33 47 53
rect 49 33 51 53
rect 69 33 71 53
rect 73 33 81 53
rect 83 33 85 53
rect 89 33 91 53
rect 93 33 101 53
rect 103 33 105 53
rect 117 33 119 53
rect 121 33 123 53
rect -19 -11 -17 9
rect -15 -11 -7 9
rect -5 -11 -3 9
rect 9 -11 11 9
rect 13 -11 15 9
rect -331 -58 -329 -38
rect -327 -58 -325 -38
rect -307 -58 -305 -38
rect -303 -58 -295 -38
rect -293 -58 -291 -38
rect -287 -58 -285 -38
rect -283 -58 -275 -38
rect -273 -58 -271 -38
rect -259 -58 -257 -38
rect -255 -58 -253 -38
rect 50 -75 52 -55
rect 54 -75 56 -55
rect 60 -75 62 -55
rect 64 -75 66 -55
rect 78 -75 80 -55
rect 82 -75 84 -55
rect 119 -132 121 -112
rect 123 -132 131 -112
rect 133 -132 135 -112
rect 147 -132 149 -112
rect 151 -132 153 -112
rect -331 -166 -329 -146
rect -327 -166 -325 -146
rect -321 -166 -319 -146
rect -317 -166 -315 -146
rect -303 -166 -301 -146
rect -299 -166 -297 -146
rect -331 -236 -329 -216
rect -327 -236 -325 -216
rect -307 -236 -305 -216
rect -303 -236 -295 -216
rect -293 -236 -291 -216
rect -287 -236 -285 -216
rect -283 -236 -275 -216
rect -273 -236 -271 -216
rect -259 -236 -257 -216
rect -255 -236 -253 -216
rect -331 -344 -329 -324
rect -327 -344 -325 -324
rect -321 -344 -319 -324
rect -317 -344 -315 -324
rect -303 -344 -301 -324
rect -299 -344 -297 -324
<< ndcontact >>
rect -335 275 -331 285
rect -325 275 -321 285
rect -263 275 -259 285
rect -253 275 -249 285
rect -199 280 -195 290
rect -189 280 -185 290
rect -127 280 -123 290
rect -117 280 -113 290
rect -311 240 -307 250
rect -301 240 -297 250
rect -291 240 -287 250
rect -281 240 -277 250
rect -271 240 -267 250
rect -175 245 -171 255
rect -165 245 -161 255
rect -155 245 -151 255
rect -145 245 -141 255
rect -135 245 -131 255
rect -335 160 -331 170
rect -315 160 -311 170
rect -307 160 -303 170
rect -297 160 -293 170
rect -90 182 -86 192
rect -80 182 -76 192
rect -217 153 -213 163
rect -197 153 -193 163
rect -189 153 -185 163
rect -179 153 -175 163
rect -18 182 -14 192
rect -8 182 -4 192
rect -66 147 -62 157
rect -56 147 -52 157
rect -46 147 -42 157
rect -36 147 -32 157
rect -26 147 -22 157
rect -335 97 -331 107
rect -325 97 -321 107
rect -263 97 -259 107
rect -253 97 -249 107
rect -154 82 -150 92
rect -144 82 -140 92
rect -134 82 -130 92
rect -126 82 -122 92
rect -116 82 -112 92
rect -311 62 -307 72
rect -301 62 -297 72
rect -291 62 -287 72
rect -281 62 -277 72
rect -271 62 -267 72
rect -86 18 -82 28
rect -66 18 -62 28
rect -58 18 -54 28
rect -48 18 -44 28
rect 41 10 45 20
rect 51 10 55 20
rect -335 -18 -331 -8
rect -315 -18 -311 -8
rect -307 -18 -303 -8
rect -297 -18 -293 -8
rect 113 10 117 20
rect 123 10 127 20
rect 65 -25 69 -15
rect 75 -25 79 -15
rect 85 -25 89 -15
rect 95 -25 99 -15
rect 105 -25 109 -15
rect -23 -41 -19 -31
rect -13 -41 -9 -31
rect -3 -41 1 -31
rect 5 -41 9 -31
rect 15 -41 19 -31
rect -335 -81 -331 -71
rect -325 -81 -321 -71
rect -263 -81 -259 -71
rect -253 -81 -249 -71
rect 46 -105 50 -95
rect 66 -105 70 -95
rect 74 -105 78 -95
rect 84 -105 88 -95
rect -311 -116 -307 -106
rect -301 -116 -297 -106
rect -291 -116 -287 -106
rect -281 -116 -277 -106
rect -271 -116 -267 -106
rect 115 -162 119 -152
rect 125 -162 129 -152
rect 135 -162 139 -152
rect 143 -162 147 -152
rect 153 -162 157 -152
rect -335 -196 -331 -186
rect -315 -196 -311 -186
rect -307 -196 -303 -186
rect -297 -196 -293 -186
rect -335 -259 -331 -249
rect -325 -259 -321 -249
rect -263 -259 -259 -249
rect -253 -259 -249 -249
rect -311 -294 -307 -284
rect -301 -294 -297 -284
rect -291 -294 -287 -284
rect -281 -294 -277 -284
rect -271 -294 -267 -284
rect -335 -374 -331 -364
rect -315 -374 -311 -364
rect -307 -374 -303 -364
rect -297 -374 -293 -364
<< pdcontact >>
rect -335 298 -331 318
rect -325 298 -321 318
rect -311 298 -307 318
rect -291 298 -287 318
rect -271 298 -267 318
rect -263 298 -259 318
rect -253 298 -249 318
rect -199 303 -195 323
rect -189 303 -185 323
rect -175 303 -171 323
rect -155 303 -151 323
rect -135 303 -131 323
rect -127 303 -123 323
rect -117 303 -113 323
rect -335 190 -331 210
rect -325 190 -321 210
rect -315 190 -311 210
rect -307 190 -303 210
rect -297 190 -293 210
rect -90 205 -86 225
rect -80 205 -76 225
rect -66 205 -62 225
rect -46 205 -42 225
rect -26 205 -22 225
rect -18 205 -14 225
rect -8 205 -4 225
rect -217 183 -213 203
rect -207 183 -203 203
rect -197 183 -193 203
rect -189 183 -185 203
rect -179 183 -175 203
rect -335 120 -331 140
rect -325 120 -321 140
rect -311 120 -307 140
rect -291 120 -287 140
rect -271 120 -267 140
rect -263 120 -259 140
rect -253 120 -249 140
rect -154 112 -150 132
rect -134 112 -130 132
rect -126 112 -122 132
rect -116 112 -112 132
rect -86 48 -82 68
rect -76 48 -72 68
rect -66 48 -62 68
rect -58 48 -54 68
rect -48 48 -44 68
rect -335 12 -331 32
rect -325 12 -321 32
rect -315 12 -311 32
rect -307 12 -303 32
rect -297 12 -293 32
rect 41 33 45 53
rect 51 33 55 53
rect 65 33 69 53
rect 85 33 89 53
rect 105 33 109 53
rect 113 33 117 53
rect 123 33 127 53
rect -23 -11 -19 9
rect -3 -11 1 9
rect 5 -11 9 9
rect 15 -11 19 9
rect -335 -58 -331 -38
rect -325 -58 -321 -38
rect -311 -58 -307 -38
rect -291 -58 -287 -38
rect -271 -58 -267 -38
rect -263 -58 -259 -38
rect -253 -58 -249 -38
rect 46 -75 50 -55
rect 56 -75 60 -55
rect 66 -75 70 -55
rect 74 -75 78 -55
rect 84 -75 88 -55
rect 115 -132 119 -112
rect 135 -132 139 -112
rect 143 -132 147 -112
rect 153 -132 157 -112
rect -335 -166 -331 -146
rect -325 -166 -321 -146
rect -315 -166 -311 -146
rect -307 -166 -303 -146
rect -297 -166 -293 -146
rect -335 -236 -331 -216
rect -325 -236 -321 -216
rect -311 -236 -307 -216
rect -291 -236 -287 -216
rect -271 -236 -267 -216
rect -263 -236 -259 -216
rect -253 -236 -249 -216
rect -335 -344 -331 -324
rect -325 -344 -321 -324
rect -315 -344 -311 -324
rect -307 -344 -303 -324
rect -297 -344 -293 -324
<< polysilicon >>
rect -193 323 -191 326
rect -169 323 -167 326
rect -159 323 -157 326
rect -149 323 -147 326
rect -139 323 -137 326
rect -121 323 -119 326
rect -329 318 -327 321
rect -305 318 -303 321
rect -295 318 -293 321
rect -285 318 -283 321
rect -275 318 -273 321
rect -257 318 -255 321
rect -329 285 -327 298
rect -329 272 -327 275
rect -305 250 -303 298
rect -295 250 -293 298
rect -285 250 -283 298
rect -275 250 -273 298
rect -257 285 -255 298
rect -193 290 -191 303
rect -193 277 -191 280
rect -257 272 -255 275
rect -169 255 -167 303
rect -159 255 -157 303
rect -149 255 -147 303
rect -139 255 -137 303
rect -121 290 -119 303
rect -121 277 -119 280
rect -169 242 -167 245
rect -159 242 -157 245
rect -149 242 -147 245
rect -139 242 -137 245
rect -305 237 -303 240
rect -295 237 -293 240
rect -285 237 -283 240
rect -275 237 -273 240
rect -84 225 -82 228
rect -60 225 -58 228
rect -50 225 -48 228
rect -40 225 -38 228
rect -30 225 -28 228
rect -12 225 -10 228
rect -329 210 -327 213
rect -319 210 -317 213
rect -301 210 -299 213
rect -211 203 -209 206
rect -201 203 -199 206
rect -183 203 -181 206
rect -329 170 -327 190
rect -319 170 -317 190
rect -301 170 -299 190
rect -84 192 -82 205
rect -211 163 -209 183
rect -201 163 -199 183
rect -183 163 -181 183
rect -84 179 -82 182
rect -329 157 -327 160
rect -319 157 -317 160
rect -301 157 -299 160
rect -60 157 -58 205
rect -50 157 -48 205
rect -40 157 -38 205
rect -30 157 -28 205
rect -12 192 -10 205
rect -12 179 -10 182
rect -211 150 -209 153
rect -201 150 -199 153
rect -183 150 -181 153
rect -60 144 -58 147
rect -50 144 -48 147
rect -40 144 -38 147
rect -30 144 -28 147
rect -329 140 -327 143
rect -305 140 -303 143
rect -295 140 -293 143
rect -285 140 -283 143
rect -275 140 -273 143
rect -257 140 -255 143
rect -148 132 -146 135
rect -138 132 -136 135
rect -120 132 -118 135
rect -329 107 -327 120
rect -329 94 -327 97
rect -305 72 -303 120
rect -295 72 -293 120
rect -285 72 -283 120
rect -275 72 -273 120
rect -257 107 -255 120
rect -257 94 -255 97
rect -148 92 -146 112
rect -138 92 -136 112
rect -120 92 -118 112
rect -148 79 -146 82
rect -138 79 -136 82
rect -120 79 -118 82
rect -80 68 -78 71
rect -70 68 -68 71
rect -52 68 -50 71
rect -305 59 -303 62
rect -295 59 -293 62
rect -285 59 -283 62
rect -275 59 -273 62
rect 47 53 49 56
rect 71 53 73 56
rect 81 53 83 56
rect 91 53 93 56
rect 101 53 103 56
rect 119 53 121 56
rect -329 32 -327 35
rect -319 32 -317 35
rect -301 32 -299 35
rect -80 28 -78 48
rect -70 28 -68 48
rect -52 28 -50 48
rect 47 20 49 33
rect -80 15 -78 18
rect -70 15 -68 18
rect -52 15 -50 18
rect -329 -8 -327 12
rect -319 -8 -317 12
rect -301 -8 -299 12
rect -17 9 -15 12
rect -7 9 -5 12
rect 11 9 13 12
rect 47 7 49 10
rect -329 -21 -327 -18
rect -319 -21 -317 -18
rect -301 -21 -299 -18
rect -17 -31 -15 -11
rect -7 -31 -5 -11
rect 11 -31 13 -11
rect 71 -15 73 33
rect 81 -15 83 33
rect 91 -15 93 33
rect 101 -15 103 33
rect 119 20 121 33
rect 119 7 121 10
rect 71 -28 73 -25
rect 81 -28 83 -25
rect 91 -28 93 -25
rect 101 -28 103 -25
rect -329 -38 -327 -35
rect -305 -38 -303 -35
rect -295 -38 -293 -35
rect -285 -38 -283 -35
rect -275 -38 -273 -35
rect -257 -38 -255 -35
rect -17 -44 -15 -41
rect -7 -44 -5 -41
rect 11 -44 13 -41
rect 52 -55 54 -52
rect 62 -55 64 -52
rect 80 -55 82 -52
rect -329 -71 -327 -58
rect -329 -84 -327 -81
rect -305 -106 -303 -58
rect -295 -106 -293 -58
rect -285 -106 -283 -58
rect -275 -106 -273 -58
rect -257 -71 -255 -58
rect -257 -84 -255 -81
rect 52 -95 54 -75
rect 62 -95 64 -75
rect 80 -95 82 -75
rect 52 -108 54 -105
rect 62 -108 64 -105
rect 80 -108 82 -105
rect 121 -112 123 -109
rect 131 -112 133 -109
rect 149 -112 151 -109
rect -305 -119 -303 -116
rect -295 -119 -293 -116
rect -285 -119 -283 -116
rect -275 -119 -273 -116
rect -329 -146 -327 -143
rect -319 -146 -317 -143
rect -301 -146 -299 -143
rect 121 -152 123 -132
rect 131 -152 133 -132
rect 149 -152 151 -132
rect 121 -165 123 -162
rect 131 -165 133 -162
rect 149 -165 151 -162
rect -329 -186 -327 -166
rect -319 -186 -317 -166
rect -301 -186 -299 -166
rect -329 -199 -327 -196
rect -319 -199 -317 -196
rect -301 -199 -299 -196
rect -329 -216 -327 -213
rect -305 -216 -303 -213
rect -295 -216 -293 -213
rect -285 -216 -283 -213
rect -275 -216 -273 -213
rect -257 -216 -255 -213
rect -329 -249 -327 -236
rect -329 -262 -327 -259
rect -305 -284 -303 -236
rect -295 -284 -293 -236
rect -285 -284 -283 -236
rect -275 -284 -273 -236
rect -257 -249 -255 -236
rect -257 -262 -255 -259
rect -305 -297 -303 -294
rect -295 -297 -293 -294
rect -285 -297 -283 -294
rect -275 -297 -273 -294
rect -329 -324 -327 -321
rect -319 -324 -317 -321
rect -301 -324 -299 -321
rect -329 -364 -327 -344
rect -319 -364 -317 -344
rect -301 -364 -299 -344
rect -329 -377 -327 -374
rect -319 -377 -317 -374
rect -301 -377 -299 -374
<< polycontact >>
rect -333 288 -329 292
rect -309 256 -305 260
rect -299 288 -295 292
rect -289 267 -285 271
rect -273 285 -269 289
rect -197 293 -193 297
rect -255 288 -251 292
rect -173 261 -169 265
rect -163 293 -159 297
rect -153 272 -149 276
rect -137 290 -133 294
rect -119 293 -115 297
rect -333 180 -329 184
rect -323 173 -319 177
rect -305 173 -301 177
rect -88 195 -84 199
rect -215 173 -211 177
rect -205 166 -201 170
rect -187 166 -183 170
rect -64 163 -60 167
rect -54 195 -50 199
rect -44 174 -40 178
rect -28 192 -24 196
rect -10 195 -6 199
rect -333 110 -329 114
rect -309 78 -305 82
rect -299 110 -295 114
rect -289 89 -285 93
rect -273 107 -269 111
rect -255 110 -251 114
rect -152 95 -148 99
rect -142 102 -138 106
rect -124 95 -120 99
rect -84 38 -80 42
rect -74 31 -70 35
rect -56 31 -52 35
rect 43 23 47 27
rect -333 2 -329 6
rect -323 -5 -319 -1
rect -305 -5 -301 -1
rect 67 -9 71 -5
rect -21 -28 -17 -24
rect -11 -21 -7 -17
rect 7 -28 11 -24
rect 77 23 81 27
rect 87 2 91 6
rect 103 20 107 24
rect 121 23 125 27
rect -333 -68 -329 -64
rect -309 -100 -305 -96
rect -299 -68 -295 -64
rect -289 -89 -285 -85
rect -273 -71 -269 -67
rect -255 -68 -251 -64
rect 48 -85 52 -81
rect 58 -92 62 -88
rect 76 -92 80 -88
rect 117 -149 121 -145
rect 127 -142 131 -138
rect 145 -149 149 -145
rect -333 -176 -329 -172
rect -323 -183 -319 -179
rect -305 -183 -301 -179
rect -333 -246 -329 -242
rect -309 -278 -305 -274
rect -299 -246 -295 -242
rect -289 -267 -285 -263
rect -273 -249 -269 -245
rect -255 -246 -251 -242
rect -333 -354 -329 -350
rect -323 -361 -319 -357
rect -305 -361 -301 -357
<< metal1 >>
rect -341 321 -243 325
rect -335 318 -331 321
rect -311 318 -307 321
rect -271 318 -267 321
rect -253 318 -249 321
rect -325 292 -321 298
rect -291 292 -287 298
rect -359 288 -333 292
rect -325 288 -299 292
rect -291 288 -277 292
rect -263 289 -259 298
rect -355 177 -351 288
rect -341 266 -338 288
rect -325 285 -321 288
rect -335 272 -331 275
rect -335 269 -321 272
rect -312 267 -289 271
rect -312 266 -308 267
rect -341 263 -308 266
rect -281 264 -277 288
rect -269 285 -259 289
rect -251 288 -243 292
rect -253 272 -249 275
rect -262 268 -249 272
rect -301 260 -258 264
rect -343 256 -309 260
rect -348 184 -344 255
rect -322 223 -319 256
rect -301 250 -297 260
rect -291 253 -267 257
rect -291 250 -287 253
rect -271 250 -267 253
rect -311 237 -307 240
rect -291 237 -287 240
rect -311 233 -287 237
rect -281 230 -277 240
rect -313 226 -266 230
rect -246 223 -243 288
rect -238 280 -235 336
rect -205 326 -107 330
rect -199 323 -195 326
rect -175 323 -171 326
rect -135 323 -131 326
rect -117 323 -113 326
rect -189 297 -185 303
rect -155 297 -151 303
rect -212 293 -197 297
rect -189 293 -163 297
rect -155 293 -141 297
rect -127 294 -123 303
rect -212 271 -209 293
rect -322 220 -243 223
rect -234 268 -209 271
rect -205 271 -202 293
rect -189 290 -185 293
rect -199 277 -195 280
rect -199 274 -185 277
rect -176 272 -153 276
rect -176 271 -172 272
rect -205 268 -172 271
rect -145 269 -141 293
rect -133 290 -123 294
rect -115 293 -107 297
rect -117 277 -113 280
rect -126 273 -113 277
rect -341 213 -287 217
rect -335 210 -331 213
rect -315 210 -311 213
rect -307 210 -303 213
rect -325 184 -321 190
rect -348 180 -333 184
rect -325 180 -311 184
rect -315 177 -311 180
rect -297 177 -293 190
rect -234 177 -231 268
rect -165 265 -122 269
rect -228 261 -173 265
rect -228 190 -225 261
rect -186 228 -183 261
rect -165 255 -161 265
rect -155 258 -131 262
rect -155 255 -151 258
rect -135 255 -131 258
rect -175 242 -171 245
rect -155 242 -151 245
rect -175 238 -151 242
rect -145 235 -141 245
rect -177 231 -130 235
rect -110 228 -107 293
rect -96 228 2 232
rect -186 225 -107 228
rect -90 225 -86 228
rect -66 225 -62 228
rect -26 225 -22 228
rect -8 225 -4 228
rect -222 206 -169 210
rect -217 203 -213 206
rect -197 203 -193 206
rect -189 203 -185 206
rect -80 199 -76 205
rect -46 199 -42 205
rect -207 177 -203 183
rect -355 173 -323 177
rect -315 173 -305 177
rect -297 173 -215 177
rect -207 173 -193 177
rect -315 170 -311 173
rect -297 170 -293 173
rect -197 170 -193 173
rect -179 170 -175 183
rect -103 195 -88 199
rect -80 195 -54 199
rect -46 195 -32 199
rect -18 196 -14 205
rect -236 165 -230 170
rect -224 166 -205 170
rect -197 166 -187 170
rect -179 166 -163 170
rect -335 157 -331 160
rect -307 157 -303 160
rect -341 153 -287 157
rect -341 143 -243 147
rect -335 140 -331 143
rect -311 140 -307 143
rect -271 140 -267 143
rect -253 140 -249 143
rect -325 114 -321 120
rect -291 114 -287 120
rect -359 110 -333 114
rect -325 110 -299 114
rect -291 110 -277 114
rect -263 111 -259 120
rect -355 -1 -351 110
rect -341 88 -338 110
rect -325 107 -321 110
rect -335 94 -331 97
rect -335 91 -321 94
rect -312 89 -289 93
rect -312 88 -308 89
rect -341 85 -308 88
rect -281 86 -277 110
rect -269 107 -259 111
rect -251 110 -243 114
rect -253 94 -249 97
rect -262 90 -249 94
rect -301 82 -258 86
rect -343 78 -309 82
rect -348 6 -344 77
rect -322 45 -319 78
rect -301 72 -297 82
rect -291 75 -267 79
rect -291 72 -287 75
rect -271 72 -267 75
rect -311 59 -307 62
rect -291 59 -287 62
rect -311 55 -287 59
rect -281 52 -277 62
rect -313 48 -266 52
rect -246 45 -243 110
rect -236 87 -233 165
rect -197 163 -193 166
rect -179 163 -175 166
rect -217 150 -213 153
rect -189 150 -185 153
rect -223 146 -169 150
rect -166 106 -163 166
rect -160 135 -106 139
rect -154 132 -150 135
rect -126 132 -122 135
rect -166 102 -142 106
rect -134 99 -130 112
rect -116 99 -112 112
rect -103 99 -100 195
rect -96 173 -93 195
rect -80 192 -76 195
rect -90 179 -86 182
rect -90 176 -76 179
rect -67 174 -44 178
rect -67 173 -63 174
rect -96 170 -63 173
rect -36 171 -32 195
rect -24 192 -14 196
rect -6 195 2 199
rect -8 179 -4 182
rect -17 175 -4 179
rect -56 167 -13 171
rect -218 95 -152 99
rect -144 95 -124 99
rect -116 95 -100 99
rect -322 42 -243 45
rect -341 35 -287 39
rect -335 32 -331 35
rect -315 32 -311 35
rect -307 32 -303 35
rect -325 6 -321 12
rect -348 2 -333 6
rect -325 2 -311 6
rect -315 -1 -311 2
rect -297 -1 -293 12
rect -218 -1 -214 95
rect -144 92 -140 95
rect -116 92 -112 95
rect -154 79 -150 82
rect -134 79 -130 82
rect -126 79 -122 82
rect -157 75 -106 79
rect -103 42 -100 95
rect -97 163 -64 167
rect -97 55 -94 163
rect -77 130 -74 163
rect -56 157 -52 167
rect -46 160 -22 164
rect -46 157 -42 160
rect -26 157 -22 160
rect -66 144 -62 147
rect -46 144 -42 147
rect -66 140 -42 144
rect -36 137 -32 147
rect -68 133 -21 137
rect -1 130 2 195
rect -77 127 2 130
rect -91 71 -38 75
rect -86 68 -82 71
rect -66 68 -62 71
rect -58 68 -54 71
rect 35 56 133 60
rect -76 42 -72 48
rect -103 38 -84 42
rect -76 38 -62 42
rect -66 35 -62 38
rect -48 35 -44 48
rect 41 53 45 56
rect 65 53 69 56
rect 105 53 109 56
rect 123 53 127 56
rect -355 -5 -323 -1
rect -315 -5 -305 -1
rect -297 -5 -214 -1
rect -155 31 -99 35
rect -315 -8 -311 -5
rect -297 -8 -293 -5
rect -335 -21 -331 -18
rect -307 -21 -303 -18
rect -341 -25 -282 -21
rect -341 -35 -243 -31
rect -335 -38 -331 -35
rect -311 -38 -307 -35
rect -271 -38 -267 -35
rect -253 -38 -249 -35
rect -325 -64 -321 -58
rect -291 -64 -287 -58
rect -359 -68 -333 -64
rect -325 -68 -299 -64
rect -291 -68 -277 -64
rect -263 -67 -259 -58
rect -355 -179 -351 -68
rect -341 -90 -338 -68
rect -325 -71 -321 -68
rect -335 -84 -331 -81
rect -335 -87 -321 -84
rect -312 -89 -289 -85
rect -312 -90 -308 -89
rect -341 -93 -308 -90
rect -281 -92 -277 -68
rect -269 -71 -259 -67
rect -251 -68 -243 -64
rect -253 -84 -249 -81
rect -262 -88 -249 -84
rect -301 -96 -258 -92
rect -343 -100 -309 -96
rect -348 -172 -344 -101
rect -322 -133 -319 -100
rect -301 -106 -297 -96
rect -291 -103 -267 -99
rect -291 -106 -287 -103
rect -271 -106 -267 -103
rect -311 -119 -307 -116
rect -291 -119 -287 -116
rect -311 -123 -287 -119
rect -281 -126 -277 -116
rect -313 -130 -266 -126
rect -246 -133 -243 -68
rect -155 -91 -152 31
rect -93 31 -74 35
rect -66 31 -56 35
rect -48 31 -32 35
rect -66 28 -62 31
rect -48 28 -44 31
rect -86 15 -82 18
rect -58 15 -54 18
rect -92 11 -38 15
rect -35 -17 -32 31
rect 51 27 55 33
rect 85 27 89 33
rect 28 23 43 27
rect 51 23 77 27
rect 85 23 99 27
rect 113 24 117 33
rect -29 12 25 16
rect -23 9 -19 12
rect 5 9 9 12
rect -35 -21 -11 -17
rect -3 -24 1 -11
rect 15 -24 19 -11
rect 28 -24 31 23
rect 35 1 38 23
rect 51 20 55 23
rect 41 7 45 10
rect 41 4 55 7
rect 64 2 87 6
rect 64 1 68 2
rect 35 -2 68 1
rect 95 -1 99 23
rect 107 20 117 24
rect 125 23 133 27
rect 123 7 127 10
rect 114 3 127 7
rect 75 -5 118 -1
rect -235 -94 -152 -91
rect -80 -28 -21 -24
rect -13 -28 7 -24
rect 15 -28 31 -24
rect -322 -136 -243 -133
rect -341 -143 -287 -139
rect -335 -146 -331 -143
rect -315 -146 -311 -143
rect -307 -146 -303 -143
rect -325 -172 -321 -166
rect -348 -176 -333 -172
rect -325 -176 -311 -172
rect -315 -179 -311 -176
rect -297 -179 -293 -166
rect -80 -179 -76 -28
rect -13 -31 -9 -28
rect 15 -31 19 -28
rect -23 -44 -19 -41
rect -3 -44 1 -41
rect 5 -44 9 -41
rect -29 -48 25 -44
rect 28 -81 31 -28
rect 34 -9 67 -5
rect 34 -69 37 -9
rect 54 -42 57 -9
rect 75 -15 79 -5
rect 85 -12 109 -8
rect 85 -15 89 -12
rect 105 -15 109 -12
rect 65 -28 69 -25
rect 85 -28 89 -25
rect 65 -32 89 -28
rect 95 -35 99 -25
rect 63 -39 110 -35
rect 130 -42 133 23
rect 54 -45 133 -42
rect 40 -52 94 -48
rect 46 -55 50 -52
rect 66 -55 70 -52
rect 74 -55 78 -52
rect 56 -81 60 -75
rect 28 -85 48 -81
rect 56 -85 70 -81
rect 66 -88 70 -85
rect 84 -88 88 -75
rect -355 -183 -323 -179
rect -315 -183 -305 -179
rect -297 -183 -76 -179
rect -5 -92 34 -88
rect -315 -186 -311 -183
rect -297 -186 -293 -183
rect -335 -199 -331 -196
rect -307 -199 -303 -196
rect -341 -203 -282 -199
rect -341 -213 -243 -209
rect -335 -216 -331 -213
rect -311 -216 -307 -213
rect -271 -216 -267 -213
rect -253 -216 -249 -213
rect -325 -242 -321 -236
rect -291 -242 -287 -236
rect -359 -246 -333 -242
rect -325 -246 -299 -242
rect -291 -246 -277 -242
rect -263 -245 -259 -236
rect -355 -357 -351 -246
rect -341 -268 -338 -246
rect -325 -249 -321 -246
rect -335 -262 -331 -259
rect -335 -265 -321 -262
rect -312 -267 -289 -263
rect -312 -268 -308 -267
rect -341 -271 -308 -268
rect -281 -270 -277 -246
rect -269 -249 -259 -245
rect -251 -246 -243 -242
rect -253 -262 -249 -259
rect -262 -266 -249 -262
rect -301 -274 -258 -270
rect -343 -278 -309 -274
rect -348 -350 -344 -279
rect -322 -311 -319 -278
rect -301 -284 -297 -274
rect -291 -281 -267 -277
rect -291 -284 -287 -281
rect -271 -284 -267 -281
rect -311 -297 -307 -294
rect -291 -297 -287 -294
rect -311 -301 -287 -297
rect -281 -304 -277 -294
rect -313 -308 -266 -304
rect -246 -311 -243 -246
rect -5 -270 -2 -92
rect 39 -92 58 -88
rect 66 -92 76 -88
rect 84 -92 106 -88
rect 66 -95 70 -92
rect 84 -95 88 -92
rect 46 -108 50 -105
rect 74 -108 78 -105
rect 40 -112 94 -108
rect 103 -138 106 -92
rect 109 -109 163 -105
rect 115 -112 119 -109
rect 143 -112 147 -109
rect 103 -142 127 -138
rect 135 -145 139 -132
rect 153 -145 157 -132
rect -233 -273 -2 -270
rect 62 -149 117 -145
rect 125 -149 145 -145
rect 153 -149 166 -145
rect -322 -314 -243 -311
rect -341 -321 -287 -317
rect -335 -324 -331 -321
rect -315 -324 -311 -321
rect -307 -324 -303 -321
rect -325 -350 -321 -344
rect -348 -354 -333 -350
rect -325 -354 -311 -350
rect -315 -357 -311 -354
rect -297 -357 -293 -344
rect 62 -357 65 -149
rect 125 -152 129 -149
rect 153 -152 157 -149
rect 115 -165 119 -162
rect 135 -165 139 -162
rect 143 -165 147 -162
rect 109 -169 163 -165
rect -355 -361 -323 -357
rect -315 -361 -305 -357
rect -297 -361 65 -357
rect -315 -364 -311 -361
rect -297 -364 -293 -361
rect -335 -377 -331 -374
rect -307 -377 -303 -374
rect -341 -381 -282 -377
<< m2contact >>
rect -348 255 -343 260
rect -258 259 -252 265
rect -240 275 -235 280
rect -122 264 -116 270
rect -228 185 -223 190
rect -230 165 -224 170
rect -348 77 -343 82
rect -258 81 -252 87
rect -236 82 -231 87
rect -13 166 -7 172
rect -97 50 -92 55
rect -348 -101 -343 -96
rect -258 -97 -252 -91
rect -99 30 -93 35
rect -240 -96 -235 -91
rect 118 -6 124 0
rect 34 -74 39 -69
rect -348 -279 -343 -274
rect -258 -275 -252 -269
rect -238 -275 -233 -269
rect 34 -93 39 -88
<< metal2 >>
rect -362 256 -348 260
rect -240 264 -235 275
rect -116 265 -102 269
rect -252 260 -235 264
rect -228 170 -224 185
rect -7 167 10 171
rect -359 78 -348 82
rect -252 82 -236 86
rect -97 35 -93 50
rect 134 49 142 53
rect 124 -5 137 -1
rect 35 -88 39 -74
rect -359 -100 -348 -96
rect -252 -96 -240 -92
rect -359 -278 -348 -274
rect -252 -274 -238 -270
<< labels >>
rlabel metal1 -292 -308 -287 -304 1 gnd
rlabel metal1 -292 -130 -287 -126 1 gnd
rlabel metal1 -292 48 -287 52 1 gnd
rlabel metal1 -292 226 -287 230 1 gnd
rlabel metal1 -330 -265 -327 -262 1 gnd
rlabel metal1 -330 -87 -327 -84 1 gnd
rlabel metal1 -330 91 -327 94 1 gnd
rlabel metal1 -259 -265 -256 -262 1 gnd
rlabel metal1 -259 -87 -256 -84 1 gnd
rlabel metal1 -259 91 -256 94 1 gnd
rlabel metal1 -259 269 -256 272 1 gnd
rlabel metal1 -317 -213 -313 -209 4 vdd
rlabel metal1 -317 -35 -313 -31 4 vdd
rlabel metal1 -317 143 -313 147 4 vdd
rlabel metal1 -317 321 -313 325 4 vdd
rlabel metal1 -341 -321 -337 -317 4 vdd
rlabel metal1 -341 -143 -337 -139 4 vdd
rlabel metal1 -341 35 -337 39 4 vdd
rlabel metal1 -341 -381 -337 -377 2 gnd
rlabel metal1 -341 -203 -337 -199 2 gnd
rlabel metal1 -341 -25 -337 -21 2 gnd
rlabel metal1 -341 213 -337 217 4 vdd
rlabel metal1 -341 153 -337 157 2 gnd
rlabel metal2 -251 82 -247 86 1 p2
rlabel metal1 -284 173 -280 177 1 g1
rlabel metal1 -359 288 -355 292 3 a1
rlabel metal1 -282 -5 -276 -1 1 g2
rlabel metal1 -157 75 -153 79 2 gnd
rlabel metal1 -159 135 -155 139 4 vdd
rlabel metal1 -156 231 -151 235 1 gnd
rlabel metal1 -194 274 -191 277 1 gnd
rlabel metal1 -123 274 -120 277 1 gnd
rlabel metal1 -181 326 -177 330 4 vdd
rlabel metal2 -105 265 -102 269 1 sum2
rlabel metal1 -223 146 -219 150 2 gnd
rlabel metal1 -222 206 -214 210 1 vdd
rlabel metal1 -86 11 -82 15 2 gnd
rlabel metal1 -91 71 -83 75 1 vdd
rlabel metal2 -252 -96 -248 -92 1 p3
rlabel metal1 -288 -183 -284 -179 1 g3
rlabel metal2 -250 -274 -246 -270 1 p4
rlabel metal1 -287 -361 -283 -357 1 g4
rlabel metal1 -47 133 -42 137 1 gnd
rlabel metal1 -85 176 -82 179 1 gnd
rlabel metal1 -14 176 -11 179 1 gnd
rlabel metal1 -72 228 -68 232 4 vdd
rlabel metal1 -28 12 -24 16 4 vdd
rlabel metal1 -26 -48 -22 -44 2 gnd
rlabel metal2 137 49 141 53 1 sum3
rlabel metal1 59 56 63 60 4 vdd
rlabel metal1 117 4 120 7 1 gnd
rlabel metal1 46 4 49 7 1 gnd
rlabel metal1 84 -39 89 -35 1 gnd
rlabel metal1 40 -112 44 -108 2 gnd
rlabel metal1 40 -52 44 -48 4 vdd
rlabel metal2 3 167 10 171 1 sum3
rlabel metal2 133 -5 137 -1 1 sum4
rlabel metal1 110 -109 114 -105 4 vdd
rlabel metal1 112 -169 116 -165 2 gnd
rlabel metal1 163 -149 166 -145 7 c5
rlabel metal1 -359 -246 -356 -242 3 a4
rlabel metal2 -359 -100 -356 -96 3 b3
rlabel metal1 -359 -68 -356 -64 3 a3
rlabel metal2 -359 78 -356 82 3 b2
rlabel metal1 -359 110 -356 114 3 a2
rlabel metal2 -359 -278 -356 -274 3 b4
rlabel metal1 -238 332 -235 336 5 sum1
rlabel metal1 -330 269 -326 272 1 gnd
rlabel metal2 -362 256 -356 260 3 b1
<< end >>
