magic
tech scmos
timestamp 1619529655
<< nwell >>
rect -184 95 -158 127
rect -141 95 -105 127
rect -93 95 -57 127
rect 18 95 54 127
rect 66 95 102 127
rect -176 21 -150 53
rect -141 21 -105 53
rect -93 21 -57 53
rect -17 21 9 53
rect 18 21 54 53
rect 66 21 102 53
<< ntransistor >>
rect -172 71 -170 81
rect -129 71 -127 81
rect -119 71 -117 81
rect -81 71 -79 81
rect -71 71 -69 81
rect 30 71 32 81
rect 40 71 42 81
rect 78 71 80 81
rect 88 71 90 81
rect -164 -3 -162 7
rect -129 -3 -127 7
rect -119 -3 -117 7
rect -81 -3 -79 7
rect -71 -3 -69 7
rect -5 -3 -3 7
rect 30 -3 32 7
rect 40 -3 42 7
rect 78 -3 80 7
rect 88 -3 90 7
<< ptransistor >>
rect -172 101 -170 121
rect -129 101 -127 121
rect -119 101 -117 121
rect -81 101 -79 121
rect -71 101 -69 121
rect 30 101 32 121
rect 40 101 42 121
rect 78 101 80 121
rect 88 101 90 121
rect -164 27 -162 47
rect -129 27 -127 47
rect -119 27 -117 47
rect -81 27 -79 47
rect -71 27 -69 47
rect -5 27 -3 47
rect 30 27 32 47
rect 40 27 42 47
rect 78 27 80 47
rect 88 27 90 47
<< ndiffusion >>
rect -174 71 -172 81
rect -170 71 -168 81
rect -131 71 -129 81
rect -127 71 -119 81
rect -117 71 -115 81
rect -83 71 -81 81
rect -79 71 -71 81
rect -69 71 -67 81
rect 28 71 30 81
rect 32 71 40 81
rect 42 71 44 81
rect 76 71 78 81
rect 80 71 88 81
rect 90 71 92 81
rect -166 -3 -164 7
rect -162 -3 -160 7
rect -131 -3 -129 7
rect -127 -3 -119 7
rect -117 -3 -115 7
rect -83 -3 -81 7
rect -79 -3 -71 7
rect -69 -3 -67 7
rect -7 -3 -5 7
rect -3 -3 -1 7
rect 28 -3 30 7
rect 32 -3 40 7
rect 42 -3 44 7
rect 76 -3 78 7
rect 80 -3 88 7
rect 90 -3 92 7
<< pdiffusion >>
rect -174 101 -172 121
rect -170 101 -168 121
rect -131 101 -129 121
rect -127 101 -125 121
rect -121 101 -119 121
rect -117 101 -115 121
rect -83 101 -81 121
rect -79 101 -77 121
rect -73 101 -71 121
rect -69 101 -67 121
rect 28 101 30 121
rect 32 101 34 121
rect 38 101 40 121
rect 42 101 44 121
rect 76 101 78 121
rect 80 101 82 121
rect 86 101 88 121
rect 90 101 92 121
rect -166 27 -164 47
rect -162 27 -160 47
rect -131 27 -129 47
rect -127 27 -125 47
rect -121 27 -119 47
rect -117 27 -115 47
rect -83 27 -81 47
rect -79 27 -77 47
rect -73 27 -71 47
rect -69 27 -67 47
rect -7 27 -5 47
rect -3 27 -1 47
rect 28 27 30 47
rect 32 27 34 47
rect 38 27 40 47
rect 42 27 44 47
rect 76 27 78 47
rect 80 27 82 47
rect 86 27 88 47
rect 90 27 92 47
<< ndcontact >>
rect -178 71 -174 81
rect -168 71 -164 81
rect -135 71 -131 81
rect -115 71 -111 81
rect -87 71 -83 81
rect -67 71 -63 81
rect 24 71 28 81
rect 44 71 48 81
rect 72 71 76 81
rect 92 71 96 81
rect -170 -3 -166 7
rect -160 -3 -156 7
rect -135 -3 -131 7
rect -115 -3 -111 7
rect -87 -3 -83 7
rect -67 -3 -63 7
rect -11 -3 -7 7
rect -1 -3 3 7
rect 24 -3 28 7
rect 44 -3 48 7
rect 72 -3 76 7
rect 92 -3 96 7
<< pdcontact >>
rect -178 101 -174 121
rect -168 101 -164 121
rect -135 101 -131 121
rect -125 101 -121 121
rect -115 101 -111 121
rect -87 101 -83 121
rect -77 101 -73 121
rect -67 101 -63 121
rect 24 101 28 121
rect 34 101 38 121
rect 44 101 48 121
rect 72 101 76 121
rect 82 101 86 121
rect 92 101 96 121
rect -170 27 -166 47
rect -160 27 -156 47
rect -135 27 -131 47
rect -125 27 -121 47
rect -115 27 -111 47
rect -87 27 -83 47
rect -77 27 -73 47
rect -67 27 -63 47
rect -11 27 -7 47
rect -1 27 3 47
rect 24 27 28 47
rect 34 27 38 47
rect 44 27 48 47
rect 72 27 76 47
rect 82 27 86 47
rect 92 27 96 47
<< polysilicon >>
rect -172 121 -170 124
rect -129 121 -127 124
rect -119 121 -117 124
rect -81 121 -79 124
rect -71 121 -69 124
rect 30 121 32 124
rect 40 121 42 124
rect 78 121 80 124
rect 88 121 90 124
rect -172 81 -170 101
rect -129 81 -127 101
rect -119 81 -117 101
rect -81 81 -79 101
rect -71 81 -69 101
rect 30 81 32 101
rect 40 81 42 101
rect 78 81 80 101
rect 88 81 90 101
rect -172 68 -170 71
rect -129 68 -127 71
rect -119 68 -117 71
rect -81 68 -79 71
rect -71 68 -69 71
rect 30 68 32 71
rect 40 68 42 71
rect 78 68 80 71
rect 88 68 90 71
rect -164 47 -162 50
rect -129 47 -127 50
rect -119 47 -117 50
rect -81 47 -79 50
rect -71 47 -69 50
rect -5 47 -3 50
rect 30 47 32 50
rect 40 47 42 50
rect 78 47 80 50
rect 88 47 90 50
rect -164 7 -162 27
rect -129 7 -127 27
rect -119 7 -117 27
rect -81 7 -79 27
rect -71 7 -69 27
rect -5 7 -3 27
rect 30 7 32 27
rect 40 7 42 27
rect 78 7 80 27
rect 88 7 90 27
rect -164 -6 -162 -3
rect -129 -6 -127 -3
rect -119 -6 -117 -3
rect -81 -6 -79 -3
rect -71 -6 -69 -3
rect -5 -6 -3 -3
rect 30 -6 32 -3
rect 40 -6 42 -3
rect 78 -6 80 -3
rect 88 -6 90 -3
<< polycontact >>
rect -176 84 -172 88
rect -133 91 -129 95
rect -123 84 -119 88
rect -85 91 -81 95
rect -75 84 -71 88
rect 26 91 30 95
rect 36 84 40 88
rect 74 91 78 95
rect 84 84 88 88
rect -168 12 -164 16
rect -133 17 -129 21
rect -123 10 -119 14
rect -85 17 -81 21
rect -75 10 -71 14
rect -9 12 -5 16
rect 26 17 30 21
rect 36 10 40 14
rect 74 17 78 21
rect 84 10 88 14
<< metal1 >>
rect -190 131 5 134
rect -190 88 -187 131
rect -184 124 -158 128
rect -141 124 -105 128
rect -93 124 -57 128
rect -178 121 -174 124
rect -135 121 -131 124
rect -115 121 -111 124
rect -87 121 -83 124
rect -67 121 -63 124
rect 2 105 5 131
rect 18 124 54 128
rect 66 124 102 128
rect 24 121 28 124
rect 44 121 48 124
rect -168 88 -164 101
rect -125 95 -121 101
rect -153 91 -133 95
rect -125 91 -111 95
rect -77 95 -73 101
rect 72 121 76 124
rect 92 121 96 124
rect 34 95 38 101
rect -98 91 -85 95
rect -77 91 -63 95
rect -194 84 -176 88
rect -168 84 -161 88
rect -168 81 -164 84
rect -178 68 -174 71
rect -184 64 -158 68
rect -153 61 -150 91
rect -115 88 -111 91
rect -67 88 -63 91
rect -23 91 26 95
rect 34 91 48 95
rect 82 95 86 101
rect 61 91 74 95
rect 82 91 96 95
rect -187 58 -150 61
rect -142 84 -123 88
rect -115 84 -75 88
rect -67 84 -51 88
rect -182 16 -179 58
rect -176 50 -150 54
rect -170 47 -166 50
rect -182 12 -168 16
rect -160 14 -156 27
rect -147 21 -144 83
rect -115 81 -111 84
rect -67 81 -63 84
rect -135 68 -131 71
rect -87 68 -83 71
rect -141 64 -105 68
rect -93 64 -57 68
rect -54 64 -51 84
rect -23 64 -20 91
rect 44 88 48 91
rect 92 88 96 91
rect 12 84 36 88
rect 44 84 84 88
rect 92 84 108 88
rect 12 82 15 84
rect 7 78 15 82
rect 44 81 48 84
rect 92 81 96 84
rect -54 61 -20 64
rect -99 60 -20 61
rect -99 58 -51 60
rect -141 50 -105 54
rect -135 47 -131 50
rect -115 47 -111 50
rect -125 21 -121 27
rect -99 21 -96 58
rect -93 50 -57 54
rect -87 47 -83 50
rect -67 47 -63 50
rect -77 21 -73 27
rect -147 17 -133 21
rect -125 17 -111 21
rect -99 17 -85 21
rect -77 17 -63 21
rect -115 14 -111 17
rect -67 14 -63 17
rect -54 14 -51 50
rect -160 10 -123 14
rect -115 10 -75 14
rect -67 10 -51 14
rect -23 16 -20 60
rect -17 50 9 54
rect -11 47 -7 50
rect -23 12 -9 16
rect -1 14 3 27
rect 12 21 15 78
rect 24 68 28 71
rect 72 68 76 71
rect 105 68 108 84
rect 18 64 54 68
rect 66 64 102 68
rect 105 64 115 68
rect 105 61 108 64
rect 60 58 108 61
rect 18 50 54 54
rect 24 47 28 50
rect 44 47 48 50
rect 34 21 38 27
rect 60 21 63 58
rect 66 50 102 54
rect 72 47 76 50
rect 92 47 96 50
rect 82 21 86 27
rect 12 17 26 21
rect 34 17 48 21
rect 60 17 74 21
rect 82 17 96 21
rect 44 14 48 17
rect 92 14 96 17
rect 105 14 108 50
rect -1 10 36 14
rect 44 10 84 14
rect 92 10 108 14
rect -160 7 -156 10
rect -115 7 -111 10
rect -67 7 -63 10
rect -1 7 3 10
rect 44 7 48 10
rect 92 7 96 10
rect -170 -6 -166 -3
rect -135 -6 -131 -3
rect -87 -6 -83 -3
rect -11 -6 -7 -3
rect 24 -6 28 -3
rect 72 -6 76 -3
rect -176 -10 -150 -6
rect -141 -10 -105 -6
rect -93 -10 -57 -6
rect -17 -10 9 -6
rect 18 -10 54 -6
rect 66 -10 102 -6
<< m2contact >>
rect -103 91 -98 96
rect 2 100 7 105
rect -161 83 -156 88
rect 56 91 61 96
rect -147 83 -142 88
rect 2 78 7 83
rect -54 50 -49 55
rect 105 50 110 55
<< metal2 >>
rect -156 84 -147 88
rect -102 58 -98 91
rect 2 83 6 100
rect 57 58 61 91
rect -102 55 -50 58
rect 57 55 109 58
rect -102 54 -54 55
rect 57 54 105 55
<< labels >>
rlabel metal1 -141 -10 -137 -6 2 gnd
rlabel metal1 18 -10 22 -6 2 gnd
rlabel metal1 -141 64 -137 68 2 gnd
rlabel metal1 18 64 22 68 2 gnd
rlabel metal1 -93 -10 -89 -6 2 gnd
rlabel metal1 66 -10 70 -6 2 gnd
rlabel metal1 -93 64 -89 68 2 gnd
rlabel metal1 66 64 70 68 2 gnd
rlabel metal1 -141 50 -137 54 4 vdd
rlabel metal1 18 50 22 54 4 vdd
rlabel metal1 -141 124 -137 128 4 vdd
rlabel metal1 18 124 22 128 4 vdd
rlabel metal1 -93 50 -89 54 4 vdd
rlabel metal1 66 50 70 54 4 vdd
rlabel metal1 -93 124 -89 128 4 vdd
rlabel metal1 66 124 70 128 4 vdd
rlabel metal1 -176 -10 -172 -6 2 gnd
rlabel metal1 -17 -10 -13 -6 2 gnd
rlabel metal1 -175 50 -171 54 4 vdd
rlabel metal1 -16 50 -12 54 4 vdd
rlabel metal1 -187 58 -179 61 3 d
rlabel metal1 105 64 115 68 7 q
rlabel metal1 -184 64 -180 68 2 gnd
rlabel metal1 -183 124 -179 128 4 vdd
rlabel metal1 -194 84 -190 88 3 clk
<< end >>
