magic
tech scmos
timestamp 1618766060
<< nwell >>
rect -6 -6 20 26
<< ntransistor >>
rect 6 -30 8 -20
<< ptransistor >>
rect 6 0 8 20
<< ndiffusion >>
rect 4 -30 6 -20
rect 8 -30 10 -20
<< pdiffusion >>
rect 4 0 6 20
rect 8 0 10 20
<< ndcontact >>
rect 0 -30 4 -20
rect 10 -30 14 -20
<< pdcontact >>
rect 0 0 4 20
rect 10 0 14 20
<< polysilicon >>
rect 6 20 8 23
rect 6 -20 8 0
rect 6 -33 8 -30
<< polycontact >>
rect 2 -15 6 -11
<< metal1 >>
rect -6 23 20 27
rect 0 20 4 23
rect 10 -6 14 0
rect 10 -10 20 -6
rect -6 -15 2 -11
rect 10 -20 14 -10
rect 0 -33 4 -30
rect -6 -37 20 -33
<< labels >>
rlabel metal1 16 -10 20 -6 7 out
rlabel metal1 -6 -15 -2 -11 3 in
rlabel metal1 -6 -37 -2 -33 2 gnd
rlabel metal1 -5 23 -1 27 4 vdd
<< end >>
